module srl 
(
	input  [31:0] rs,
	input  [4: 0] shamt,
	output [31:0] rd
);
assign rd = rs >> shamt;
endmodule
